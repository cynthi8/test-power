`timescale 1ns/1ps
`celldefine
module DHFILLHLHLS11();


endmodule
`endcelldefine
