`timescale 1ns/1ps
`celldefine
module CLOAD1 (INP);
input INP;



endmodule
`endcelldefine
