`timescale 1ns/1ps
`celldefine
module HEADX4 (SLEEP);
input SLEEP;



endmodule
`endcelldefine
