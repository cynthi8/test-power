`timescale 1ns/1ps
`celldefine
module HEADX8 (SLEEP);
input SLEEP;



endmodule
`endcelldefine
