`timescale 1ns/1ps
`celldefine
module TIEH (Z);
output Z;



endmodule
`endcelldefine
