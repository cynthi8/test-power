`timescale 1ns/1ps
`celldefine
module SHFILL1();


endmodule
`endcelldefine
