`timescale 1ns/1ps
`celldefine
module DCAP();


endmodule
`endcelldefine
