`timescale 1ns/1ps
`celldefine
module SHFILL64();


endmodule
`endcelldefine
