`timescale 1ns/1ps
`celldefine
module SHFILL2();


endmodule
`endcelldefine
