`timescale 1ns/1ps
`celldefine
module DHFILLHLH2();


endmodule
`endcelldefine
