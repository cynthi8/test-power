`timescale 1ns/1ps
`celldefine
module HEADX16 (SLEEP);
input SLEEP;



endmodule
`endcelldefine
