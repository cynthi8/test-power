`timescale 1ns/1ps
`celldefine
module BUSKP (INP);
input INP;



endmodule
`endcelldefine
