`timescale 1ns/1ps
`celldefine
module HEADX2 (SLEEP);
input SLEEP;



endmodule
`endcelldefine
