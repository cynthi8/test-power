`timescale 1ns/1ps
`celldefine
module NMT3 (G, D, S);
input G;
input D;
input S;



endmodule
`endcelldefine
