`timescale 1ns/1ps
`celldefine
module TIEL (ZN);
output ZN;



endmodule
`endcelldefine
