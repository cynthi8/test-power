`timescale 1ns/1ps
`celldefine
module HEADX32 (SLEEP);
input SLEEP;



endmodule
`endcelldefine
