`timescale 1ns/1ps
`celldefine
module DHFILLLHL2();


endmodule
`endcelldefine
