`timescale 1ns/1ps
`celldefine
module ANTENNA (INP);
input INP;



endmodule
`endcelldefine
