`timescale 1ns/1ps
`celldefine
module PMT1 (G, D, S);
input G;
input D;
input S;



endmodule
`endcelldefine
