`timescale 1ns/1ps
`celldefine
module SHFILL128();


endmodule
`endcelldefine
