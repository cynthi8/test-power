`timescale 1ns/1ps
`celldefine
module SHFILL3();


endmodule
`endcelldefine
